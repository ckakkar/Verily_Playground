module hello;

initial begin
    $display("Hello, Verilog on Mac!");
    $finish;
end

endmodule